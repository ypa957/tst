module compare

endmodule